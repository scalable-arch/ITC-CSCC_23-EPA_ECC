module GFMULT(a, b, c);
  input [7:0] a;
  input [7:0] b;
  output [7:0] c;

  /*
    GF(2^8)
    primitive polynomial : x^8 + x6 + x^4 + x^3 + x^2 + x + 1 => Unity ECC와 같다.
    a = a^n
    b = a^m
    c = a^(n+m)
  */

  assign c = ({8{b[0]}} & ((a << 0))) ^
  ({8{b[1]}} & ((a << 1) ^ ({8{a[7]}} & 8'b0101_1111))) ^ 
  ({8{b[2]}} & ((a << 2) ^ ({8{a[7]}} & 8'b1011_1110) ^ ({8{a[6]}} & 8'b0101_1111))) ^ 
  ({8{b[3]}} & ((a << 3) ^ ({8{a[7]}} & 8'b0010_0011) ^ ({8{a[6]}} & 8'b1011_1110) ^ ({8{a[5]}} & 8'b0101_1111))) ^
  ({8{b[4]}} & ((a << 4) ^ ({8{a[7]}} & 8'b0100_0110) ^ ({8{a[6]}} & 8'b0010_0011) ^ ({8{a[5]}} & 8'b1011_1110) ^ ({8{a[4]}} & 8'b0101_1111))) ^
  ({8{b[5]}} & ((a << 5) ^ ({8{a[7]}} & 8'b1000_1100) ^ ({8{a[6]}} & 8'b0100_0110) ^ ({8{a[5]}} & 8'b0010_0011) ^ ({8{a[4]}} & 8'b1011_1110) ^ ({8{a[3]}} & 8'b0101_1111))) ^
  ({8{b[6]}} & ((a << 6) ^ ({8{a[7]}} & 8'b0100_0111) ^ ({8{a[6]}} & 8'b1000_1100) ^ ({8{a[5]}} & 8'b0100_0110) ^ ({8{a[4]}} & 8'b0010_0011) ^ ({8{a[3]}} & 8'b1011_1110) ^ ({8{a[2]}} & 8'b0101_1111))) ^ 
  ({8{b[7]}} & ((a << 7) ^ ({8{a[7]}} & 8'b1000_1110) ^ ({8{a[6]}} & 8'b0100_0111) ^ ({8{a[5]}} & 8'b1000_1100) ^ ({8{a[4]}} & 8'b0100_0110) ^ ({8{a[3]}} & 8'b0010_0011) ^ ({8{a[2]}} & 8'b1011_1110) ^ ({8{a[1]}} & 8'b0101_1111)));
endmodule