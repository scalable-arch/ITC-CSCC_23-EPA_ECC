
module SEC_DED_ENCODER(input [95:0] data_in, output [103:0] codeword_out);

	assign codeword_out[103:8] = data_in[95:0];
	assign codeword_out[7] = ^(data_in&96'b111111111111111111111000000000000000000000000000000000001111111111111111111111111111111111100000);
	assign codeword_out[6] = ^(data_in&96'b111111000000000000000111111111111111000000000000000000001111111111111111111100000000000000011111);
	assign codeword_out[5] = ^(data_in&96'b100000111110000000000111110000000000111111111100000000001111111111000000000011111111110000011111);
	assign codeword_out[4] = ^(data_in&96'b010000100001111000000100001111000000111100000011111100001111000000111111000011111100001111011111);
	assign codeword_out[3] = ^(data_in&96'b001000010001000111000010001000111000100011100011100011101000111000111000111011100011101110111100);
	assign codeword_out[2] = ^(data_in&96'b000100001000100100110001000100100110010010011010011011010100100110100110110110011011011101110011);
	assign codeword_out[1] = ^(data_in&96'b000010000100010010101000100010010101001001010101010110110010010101010101101101010110111011101010);
	assign codeword_out[0] = ^(data_in&96'b000001000010001001011000010001001011000100101100101101110001001011001011011100101101110111100101);

endmodule


